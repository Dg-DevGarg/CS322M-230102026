`timescale 1ns/1ns
module L1_2(input [3:0] A,B,output result);
  assign result = A==B;
endmodule
